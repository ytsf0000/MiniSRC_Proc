module Register (
	input clk,
	input reset,
	input enable
	
);

endmodule