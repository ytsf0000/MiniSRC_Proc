module CLA_32B (
	input[31:0] a,
	input[31:0] b
);

endmodule