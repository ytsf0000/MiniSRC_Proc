module RegisterFile(
	input [4:0] ra,
	input [4:0] rb,
	input [4:0] rc,
	input rin,
	input rout,
	output [31:0] BusMuxOut
);

	

endmodule 