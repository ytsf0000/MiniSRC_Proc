module MIPS_Proc ();

endmodule