module ALU_Shifting (
	input [32:0] a,
	input SHR,
	input SHRA,
	input SHL,
	input ROR,
	input ROL,
	output [32:0] c
);

endmodule