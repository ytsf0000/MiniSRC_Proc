module ALU_Logical_tb ();

	reg in_and;
	reg in_or;
	reg in_neg;
	reg in_not;
	reg [31:0] a;
	reg [31:0] b;
	wire [31:0] c;

endmodule