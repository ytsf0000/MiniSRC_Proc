module AddSub_64B_tb ();

	reg [128:0] stimulus;
	reg [64:0] test_sum;
	reg clk;

	//output values
	wire signed [63:0] s; // sum
	wire signed [63:0] x;
	wire signed [63:0] y;
	wire c_out; //c4 is c_out
	wire g; // for higher-bit compound CLA 
	wire p;
	
	assign x = stimulus[63:0];
	assign y = stimulus[127:64];
	
	// It is obviously unrealistic to provide all 2^(16+16+1) arithmetic operations, so a pseudo-randomized pool of cases are chosen instead.
	// 10000 cases are generated by a 32-bit LFSR.
	
	always @ (posedge clk) begin
		stimulus <= {stimulus[31:0], stimulus[32] ^ stimulus[19] ^ stimulus[18] ^ stimulus[1]};
	end
	
	// testbench correctness assertion
	always @ (posedge clk) begin
		$display("Test case: x = %d, y = %d, c_in = %d, sum = %d, c_out = %d", x, y, stimulus[32], s, c_out);
		test_sum = {1'b0,x} + {1'b0,y} + {16'b0,stimulus[32]};
		if (!(test_sum[15:0] == s)) begin
			$display("Sum is incorrect, expected %d when given sum of %d", test_sum, s);
			$finish;
		end
		if (!(test_sum[16] == c_out)) begin
			$display("Incorrect carry signal, expected: %b, instead got: %b", test_sum[16], c_out);
			$finish;
		end
	end
	
	initial begin
		stimulus <= 33'b1;
		clk <= 1'b0;
		repeat (10000) begin
			#10;
			clk <= 1'b1;
			#10;
			clk <= 1'b0;
		end
		
		$display("Testbench complete.");
	end
	
	SixteenBitCLA test_16b_CLA(
		.x(stimulus[15:0]),
		.y(stimulus[31:16]),
		.c_in(stimulus[32]),
		.s(s), // sum
		.c_out(c_out), //c4 is c_out
		.g(g), // for higher-bit compound CLA 
		.p(p)
	);

endmodule
