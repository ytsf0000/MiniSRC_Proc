module CLA_64B_tb();

	reg [128:0] stimulus;
	reg [64:0] test_sum;
	reg clk;

	//output values
	wire signed [63:0] s; // sum
	wire signed [63:0] x;
	wire signed [63:0] y;
	wire c_out; //c4 is c_out
	
	assign x = stimulus[63:0];
	assign y = stimulus[127:64];
	
	CLA_64B test_CLA_64B(
		.a(stimulus[63:0]),
		.b(stimulus[127:64]),
		.c_in(stimulus[128]),
		.s(s), // sum
		.c_out(c_out) //c4 is c_out
	);
	
	// It is obviously unrealistic to provide all 2^(16+16+1) arithmetic operations, so a pseudo-randomized pool of cases are chosen instead.
	// 10000 cases are generated by a 32-bit LFSR.
	
	always @ (posedge clk) begin
		stimulus <= {stimulus[127:0],~(stimulus[128]^stimulus[123])};
	end
	
	// testbench correctness assertion
	always @ (posedge clk) begin
		$display("Test case: x = %d, y = %d, c_in = %d, sum = %d, c_out = %d", x, y, stimulus[128], s, c_out);
		test_sum = {1'b0,x} + {1'b0,y} + {64'b0,stimulus[128]};
		if (!(test_sum[63:0] == s)) begin
			$display("Sum is incorrect, expected %d when given sum of %d", test_sum, s);
			$finish;
		end
		if (!(test_sum[64] == c_out)) begin
			$display("Incorrect carry signal, expected: %b, instead got: %b", test_sum[64], c_out);
			$finish;
		end
	end
	
	initial begin
		stimulus <= 129'b1;
		clk <= 1'b0;
		repeat (10000) begin
			#10;
			clk <= 1'b1;
			#10;
			clk <= 1'b0;
		end
		
		$display("Testbench complete.");
	end

endmodule